# ====================================================================
#
#      btree.cdl
#
#      BTree library configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2018 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jturnsek 
# Contributors:   
# Date:           2018-07-18
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_BTREE_LIB {
    display         "BTree library"
    include_dir     cyg/db/btree

    requires        CYGPKG_POSIX
    requires        CYGPKG_ISOINFRA
    requires        CYGPKG_MEMALLOC
    requires        CYGPKG_LINUX_COMPAT
    requires        CYGPKG_ERROR
    requires        CYGPKG_FS_JFFS2
    
    compile         -library=libextras.a btree.c

    cdl_option CYGDAT_BTREE_LIB_PAGESIZE {
        display       "Size of the page"
        flavor        data
        default_value 512
        legal_values 512 1024 2048 4096

        description   "
            This option sets the size of the page."
    }

    cdl_option CYGDAT_BTREE_LIB_COMMIT_PAGES {
        display       "Number of commit pages"
        flavor        data
        default_value 16
        legal_values 8 16 32 64

        description   "
            This option sets the max number of pages to write in one commit."
    }

    cdl_option CYGDAT_BTREE_LIB_MAXCACHE {
        display       "Number of max cache pages"
        flavor        data
        default_value 16
        legal_values 8 16 32 64 128 256 512 1024

        description   "
            This option sets the max number of pages to keep in cache."
    }

}

# ====================================================================
# End of btree.cdl
